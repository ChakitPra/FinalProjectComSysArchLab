module ascii_rom (
    input [7:0] ascii_code,   // ASCII character input
    input [3:0] row,          // Row of the character pixel (0-15)
    output reg [7:0] pixels   // 8 pixels in the row (1 byte)
);

    reg [7:0] rom [0:127][0:15]; // ROM for 128 ASCII characters, each with 16 rows of 8 pixels

    initial begin

         // code x30 (0)
            rom[48][0]   = 8'b00000000; //
            rom[48][1]   = 8'b00000000; //
            rom[48][2]   = 8'b00111000; //  ***  
            rom[48][3]   = 8'b01101100; // ** **
            rom[48][4]   = 8'b11000110; //**   **
            rom[48][5]   = 8'b11000110; //**   **
            rom[48][6]   = 8'b11000110; //**   **
            rom[48][7]   = 8'b11000110; //**   **
            rom[48][8]   = 8'b11000110; //**   **
            rom[48][9]   = 8'b11000110; //**   **
            rom[48][10] = 8'b01101100;  // ** **
            rom[48][11] = 8'b00111000;  //  ***
            rom[48][12] = 8'b00000000;  //
            rom[48][13] = 8'b00000000;  //
            rom[48][14] = 8'b00000000;  //
            rom[48][15] = 8'b00000000;  //
            // code x31 (1)
            rom[49][0]   = 8'b00000000; //
            rom[49][1]   = 8'b00000000; //
            rom[49][2]   = 8'b00011000; //   **  
            rom[49][3]   = 8'b00111000; //  ***
            rom[49][4]   = 8'b01111000; // ****
            rom[49][5]   = 8'b00011000; //   **
            rom[49][6]   = 8'b00011000; //   **
            rom[49][7]   = 8'b00011000; //   **
            rom[49][8]   = 8'b00011000; //   **
            rom[49][9]   = 8'b00011000; //   **
            rom[49][10] = 8'b01111110;  // ******
            rom[49][11] = 8'b01111110;  // ******
            rom[49][12] = 8'b00000000;  //
            rom[49][13] = 8'b00000000;  //
            rom[49][14] = 8'b00000000;  //
            rom[49][15]= 8'b00000000;   //
            // code x32 (2)
            rom[50][0]   = 8'b00000000; //
            rom[50][1]   = 8'b00000000; //
            rom[50][2]   = 8'b11111110; //*******  
            rom[50][3]   = 8'b11111110; //*******
            rom[50][4]   = 8'b00000110; //     **
            rom[50][5]   = 8'b00000110; //     **
            rom[50][6]   = 8'b11111110; //*******
            rom[50][7]   = 8'b11111110; //*******
            rom[50][8]   = 8'b11000000; //**
            rom[50][9]   = 8'b11000000; //**
            rom[50][10] = 8'b11111110;  //*******
            rom[50][11] = 8'b11111110;  //*******
            rom[50][12] = 8'b00000000;  //
            rom[50][13] = 8'b00000000;  //
            rom[50][14] = 8'b00000000;  //
            rom[50][15] = 8'b00000000;  //
            // code x33 (3)
            rom[51][0]   = 8'b00000000; //
            rom[51][1]   = 8'b00000000; //
            rom[51][2]   = 8'b11111110; //*******  
            rom[51][3]   = 8'b11111110; //*******
            rom[51][4]   = 8'b00000110; //     **
            rom[51][5]   = 8'b00000110; //     **
            rom[51][6]   = 8'b00111110; //  *****
            rom[51][7]   = 8'b00111110; //  *****
            rom[51][8]   = 8'b00000110; //     **
            rom[51][9]   = 8'b00000110; //     **
            rom[51][10] = 8'b11111110;  //*******
            rom[51][11] = 8'b11111110;  //*******
            rom[51][12] = 8'b00000000;  //
            rom[51][13] = 8'b00000000;  //
            rom[51][14] = 8'b00000000;  //
            rom[51][15] = 8'b00000000;  //
            // code x34 (4)
            rom[52][0]   = 8'b00000000; //
            rom[52][1]   = 8'b00000000; //
            rom[52][2]   = 8'b11000110; //**   **  
            rom[52][3]   = 8'b11000110; //**   **
            rom[52][4]   = 8'b11000110; //**   **
            rom[52][5]   = 8'b11000110; //**   **
            rom[52][6]   = 8'b11111110; //*******
            rom[52][7]   = 8'b11111110; //*******
            rom[52][8]   = 8'b00000110; //     **
            rom[52][9]   = 8'b00000110; //     **
            rom[52][10] = 8'b00000110;  //     **
            rom[52][11] = 8'b00000110;  //     **
            rom[52][12] = 8'b00000000;  //
            rom[52][13] = 8'b00000000;  //
            rom[52][14] = 8'b00000000;  //
            rom[52][15]= 8'b00000000;   //
            // code x35 (5)
            rom[53][0]   = 8'b00000000; //
            rom[53][1]   = 8'b00000000; //
            rom[53][2]   = 8'b11111110; //*******  
            rom[53][3]   = 8'b11111110; //*******
            rom[53][4]   = 8'b11000000; //**
            rom[53][5]   = 8'b11000000; //**
            rom[53][6]   = 8'b11111110; //*******
            rom[53][7]   = 8'b11111110; //*******
            rom[53][8]   = 8'b00000110; //     **
            rom[53][9]   = 8'b00000110; //     **
            rom[53][10] = 8'b11111110;  //*******
            rom[53][11] = 8'b11111110;  //*******
            rom[53][12] = 8'b00000000;  //
            rom[53][13] = 8'b00000000;  //
            rom[53][14] = 8'b00000000;  //
            rom[53][15] = 8'b00000000;  //
            // code x36 (6)
            rom[54][0]   = 8'b00000000; //
            rom[54][1]   = 8'b00000000; //
            rom[54][2]   = 8'b11111110; //*******  
            rom[54][3]   = 8'b11111110; //*******
            rom[54][4]   = 8'b11000000; //**
            rom[54][5]   = 8'b11000000; //**
            rom[54][6]   = 8'b11111110; //*******
            rom[54][7]   = 8'b11111110; //*******
            rom[54][8]   = 8'b11000110; //**   **
            rom[54][9]   = 8'b11000110; //**   **
            rom[54][10] = 8'b11111110;  //*******
            rom[54][11] = 8'b11111110;  //*******
            rom[54][12] = 8'b00000000;  //
            rom[54][13] = 8'b00000000;  //
            rom[54][14] = 8'b00000000;  //
            rom[54][15] = 8'b00000000;  //
            // code x37 (7)
            rom[55][0]   = 8'b00000000; //
            rom[55][1]   = 8'b00000000; //
            rom[55][2]   = 8'b11111110; //*******  
            rom[55][3]   = 8'b11111110; //*******
            rom[55][4]   = 8'b00000110; //     **
            rom[55][5]   = 8'b00000110; //     **
            rom[55][6]   = 8'b00000110; //     **
            rom[55][7]   = 8'b00000110; //     **
            rom[55][8]   = 8'b00000110; //     **
            rom[55][9]   = 8'b00000110; //     **
            rom[55][10] = 8'b00000110;  //     **
            rom[55][11] = 8'b00000110;  //     **
            rom[55][12] = 8'b00000000;  //
            rom[55][13] = 8'b00000000;  //
            rom[55][14] = 8'b00000000;  //
            rom[55][15] = 8'b00000000;  //
            // code x38 (8)
            rom[56][0]   = 8'b00000000; //
            rom[56][1]   = 8'b00000000; //
            rom[56][2]   = 8'b11111110; //*******  
            rom[56][3]   = 8'b11111110; //*******
            rom[56][4]   = 8'b11000110; //**   **
            rom[56][5]   = 8'b11000110; //**   **
            rom[56][6]   = 8'b11111110; //*******
            rom[56][7]   = 8'b11111110; //*******
            rom[56][8]   = 8'b11000110; //**   **
            rom[56][9]   = 8'b11000110; //**   **
            rom[56][10] = 8'b11111110;  //*******
            rom[56][11] = 8'b11111110;  //*******
            rom[56][12] = 8'b00000000;  //
            rom[56][13] = 8'b00000000;  //
            rom[56][14] = 8'b00000000;  //
            rom[56][15]= 8'b00000000;   //
            // code x39 (9)
            rom[57][0]   = 8'b00000000; //
            rom[57][1]   = 8'b00000000; //
            rom[57][2]   = 8'b11111110; //*******  
            rom[57][3]   = 8'b11111110; //*******
            rom[57][4]   = 8'b11000110; //**   **
            rom[57][5]   = 8'b11000110; //**   **
            rom[57][6]   = 8'b11111110; //*******
            rom[57][7]   = 8'b11111110; //*******
            rom[57][8]   = 8'b00000110; //     **
            rom[57][9]   = 8'b00000110; //     **
            rom[57][10] = 8'b11111110;  //*******
            rom[57][11] = 8'b11111110;  //*******
            rom[57][12] = 8'b00000000;  //
            rom[57][13] = 8'b00000000;  //
            rom[57][14] = 8'b00000000;  //
            rom[57][15]= 8'b00000000;   //
            // code x41 (A)
            rom[65][0]   = 8'b00000000; //
            rom[65][1]   = 8'b00000000; //
            rom[65][2]   = 8'b00010000; //   *
            rom[65][3]   = 8'b00111000; //  ***
            rom[65][4]   = 8'b01101100; // ** **   
            rom[65][5]   = 8'b11000110; //**   **   
            rom[65][6]   = 8'b11000110; //**   **
            rom[65][7]   = 8'b11111110; //*******
            rom[65][8]   = 8'b11111110; //*******
            rom[65][9]   = 8'b11000110; //**   **
            rom[65][10] = 8'b11000110;  //**   **
            rom[65][11] = 8'b11000110;  //**   **
            rom[65][12] = 8'b00000000;  //
            rom[65][13] = 8'b00000000;  //
            rom[65][14] = 8'b00000000;  //
            rom[65][15]= 8'b00000000;   //
            // code x42 (B)
            rom[66][0]   = 8'b00000000; //
            rom[66][1]   = 8'b00000000; //
            rom[66][2]   = 8'b11111100; //******
            rom[66][3]   = 8'b11111110; //*******
            rom[66][4]   = 8'b11000110; //**   **
            rom[66][5]   = 8'b11000110; //**   **   
            rom[66][6]   = 8'b11111100; //******
            rom[65][7]   = 8'b11111100; //******
            rom[66][8]   = 8'b11000110; //**   **
            rom[66][9]   = 8'b11000110; //**   **
            rom[66][10] = 8'b11111110;  //*******
            rom[66][11] = 8'b11111100;  //******
            rom[66][12] = 8'b00000000;  //
            rom[66][13] = 8'b00000000;  //
            rom[66][14] = 8'b00000000;  //
            rom[66][15]= 8'b00000000;   //
            // code x43 (C)
            rom[67][0]   = 8'b00000000; //
            rom[67][1]   = 8'b00000000; //
            rom[67][2]   = 8'b01111100; // *****
            rom[67][3]   = 8'b11111110; //*******
            rom[67][4]   = 8'b11000000; //**
            rom[67][5]   = 8'b11000000; //**   
            rom[67][6]   = 8'b11000000; //**
            rom[67][7]   = 8'b11000000; //**
            rom[67][8]   = 8'b11000000; //** 
            rom[67][9]   = 8'b11000000; //** 
            rom[67][10] = 8'b11111110;  //*******
            rom[67][11] = 8'b01111100;  // *****
            rom[67][12] = 8'b00000000;  //
            rom[67][13] = 8'b00000000;  //
            rom[67][14] = 8'b00000000;  //
            rom[67][15]= 8'b00000000;   //
            // code x44 (D)
            rom[68][0]   = 8'b00000000; //
            rom[68][1]   = 8'b00000000; //
            rom[68][2]   = 8'b11111100; //******
            rom[68][3]   = 8'b11111110; //*******
            rom[68][4]   = 8'b11000110; //**   **
            rom[68][5]   = 8'b11000110; //**   **   
            rom[68][6]   = 8'b11000110; //**   **
            rom[68][7]   = 8'b11000110; //**   **
            rom[68][8]   = 8'b11000110; //**   ** 
            rom[68][9]   = 8'b11000110; //**   ** 
            rom[68][10] = 8'b11111110;  //*******
            rom[68][11] = 8'b11111100;  //******
            rom[68][12] = 8'b00000000;  //
            rom[68][13] = 8'b00000000;  //
            rom[68][14] = 8'b00000000;  //
            rom[68][15] = 8'b00000000;  //
            // code x45 (E)
            rom[69][0]   = 8'b00000000; //
            rom[69][1]   = 8'b00000000; //
            rom[69][2]   = 8'b11111110; //*******
            rom[69][3]   = 8'b11111110; //*******
            rom[69][4]   = 8'b11000000; //**
            rom[69][5]   = 8'b11000000; //**   
            rom[69][6]   = 8'b11111100; //******
            rom[69][7]   = 8'b11111100; //******
            rom[69][8]   = 8'b11000000; //** 
            rom[69][9]   = 8'b11000000; //** 
            rom[69][10] = 8'b11111110;  //*******
            rom[69][11] = 8'b11111110;  //*******
            rom[69][12] = 8'b00000000;  //
            rom[69][13] = 8'b00000000;  //
            rom[69][14] = 8'b00000000;  //
            rom[69][15] = 8'b00000000;  //
            // code x46 (F)
            rom[70][0]   = 8'b00000000; //
            rom[70][1]   = 8'b00000000; //
            rom[70][2]   = 8'b11111110; //*******
            rom[70][3]   = 8'b11111110; //*******
            rom[70][4]   = 8'b11000000; //**
            rom[70][5]   = 8'b11000000; //**   
            rom[70][6]   = 8'b11111100; //******
            rom[70][7]   = 8'b11111100; //******
            rom[70][8]   = 8'b11000000; //** 
            rom[70][9]   = 8'b11000000; //** 
            rom[70][10] = 8'b11000000;  //**
            rom[70][11] = 8'b11000000;  //**
            rom[70][12] = 8'b00000000;  //
            rom[70][13] = 8'b00000000;  //
            rom[70][14] = 8'b00000000;  //
            rom[70][15]= 8'b00000000;   //
            // code x47 (G)
            rom[71][0]   = 8'b00000000; //
            rom[71][1]   = 8'b00000000; //
            rom[71][2]   = 8'b01111100; // *****
            rom[71][3]   = 8'b11111110; //*******
            rom[71][4]   = 8'b11000000; //**
            rom[71][5]   = 8'b11000000; //**   
            rom[71][6]   = 8'b11111110; //*******
            rom[71][7]   = 8'b11111110; //*******
            rom[71][8]   = 8'b11000110; //**   **
            rom[71][9]   = 8'b11000110; //**   **
            rom[71][10] = 8'b11111110;  //*******
            rom[71][11] = 8'b01110110;  // *** **
            rom[71][12] = 8'b00000000;  //
            rom[71][13] = 8'b00000000;  //
            rom[71][14] = 8'b00000000;  //
            rom[71][15] = 8'b00000000;  //
            // code x48 (H)
            rom[72][0]   = 8'b00000000; //
            rom[72][1]   = 8'b00000000; //
            rom[72][2]   = 8'b11000110; //**   **
            rom[72][3]   = 8'b11000110; //**   **
            rom[72][4]   = 8'b11000110; //**   **
            rom[72][5]   = 8'b11000110; //**   **
            rom[72][6]   = 8'b11111110; //*******
            rom[72][7]   = 8'b11111110; //*******
            rom[72][8]   = 8'b11000110; //**   **
            rom[72][9]   = 8'b11000110; //**   **
            rom[72][10] = 8'b11000110;  //**   **
            rom[72][11] = 8'b11000110;  //**   **
            rom[72][12] = 8'b00000000;  //
            rom[72][13] = 8'b00000000;  //
            rom[72][14] = 8'b00000000;  //
            rom[72][15] = 8'b00000000;  //
            // code x49 (I)
            rom[73][0]   = 8'b00000000; //
            rom[73][1]   = 8'b00000000; //
            rom[73][2]   = 8'b11111110; //*******
            rom[73][3]   = 8'b11111110; //*******
            rom[73][4]   = 8'b00110000; //  **
            rom[73][5]   = 8'b00110000; //  **
            rom[73][6]   = 8'b00110000; //  **
            rom[73][7]   = 8'b00110000; //  **
            rom[73][8]   = 8'b00110000; //  **
            rom[73][9]   = 8'b00110000; //  **
            rom[73][10] = 8'b11111110;  //*******
            rom[73][11] = 8'b11111110;  //*******
            rom[73][12] = 8'b00000000;  //
            rom[73][13] = 8'b00000000;  //
            rom[73][14] = 8'b00000000;  //
            rom[73][15]= 8'b00000000;   //
            // code x4a (J)
            rom[74][0]   = 8'b00000000; //
            rom[74][1]   = 8'b00000000; //
            rom[74][2]   = 8'b11111110; //*******
            rom[74][3]   = 8'b11111110; //*******
            rom[74][4]   = 8'b00011000; //   **
            rom[74][5]   = 8'b00011000; //   **
            rom[74][6]   = 8'b00011000; //   **
            rom[74][7]   = 8'b00011000; //   **
            rom[74][8]   = 8'b00011000; //   **
            rom[74][9]   = 8'b00011000; //   **
            rom[74][10] = 8'b11111000;  //*****
            rom[74][11] = 8'b01111000;  // ****
            rom[74][12] = 8'b00000000;  //
            rom[74][13] = 8'b00000000;  //
            rom[74][14] = 8'b00000000;  //
            rom[74][15]= 8'b00000000;   //
            // code x4b (K)
            rom[75][0]   = 8'b00000000; //
            rom[75][1]   = 8'b00000000; //
            rom[75][2]   = 8'b11000110; //**   **
            rom[75][3]   = 8'b11001100; //**  **
            rom[75][4]   = 8'b11011000; //** **
            rom[75][5]   = 8'b11110000; //****
            rom[75][6]   = 8'b11100000; //***
            rom[75][7]   = 8'b11100000; //***
            rom[75][8]   = 8'b11110000; //****
            rom[75][9]   = 8'b11011000; //** **
            rom[75][10] = 8'b11001100;  //**  **
            rom[75][11] = 8'b11000110;  //**   **
            rom[75][12] = 8'b00000000;  //
            rom[75][13] = 8'b00000000;  //
            rom[75][14] = 8'b00000000;  //
            rom[75][15] = 8'b00000000;  //
            // code x4c (L)
            rom[76][0]   = 8'b00000000; //
            rom[76][1]   = 8'b00000000; //
            rom[76][2]   = 8'b11000000; //**
            rom[76][3]   = 8'b11000000; //**
            rom[76][4]   = 8'b11000000; //**
            rom[76][5]   = 8'b11000000; //**
            rom[76][6]   = 8'b11000000; //**
            rom[76][7]   = 8'b11000000; //**
            rom[76][8]   = 8'b11000000; //**
            rom[76][9]   = 8'b11000000; //**
            rom[76][10] = 8'b11111110;  //*******
            rom[76][11] = 8'b11111110;  //*******
            rom[76][12] = 8'b00000000;  //
            rom[76][13] = 8'b00000000;  //
            rom[76][14] = 8'b00000000;  //
            rom[76][15]= 8'b00000000;   //
            // code x4d (M)
            rom[77][0]   = 8'b00000000; //
            rom[77][1]   = 8'b00000000; //
            rom[77][2]   = 8'b11000110; //**   **
            rom[77][3]   = 8'b11000110; //**   **
            rom[77][4]   = 8'b11101110; //*** ***
            rom[77][5]   = 8'b11111110; //*******
            rom[77][6]   = 8'b11010110; //** * **
            rom[77][7]   = 8'b11000110; //**   **
            rom[77][8]   = 8'b11000110; //**   **
            rom[77][9]   = 8'b11000110; //**   **
            rom[77][10] = 8'b11000110;  //**   **
            rom[77][11] = 8'b11000110;  //**   **
            rom[77][12] = 8'b00000000;  //
            rom[77][13] = 8'b00000000;  //
            rom[77][14] = 8'b00000000;  //
            rom[77][15] = 8'b00000000;  //
            // code x4e (N)
            rom[78][0]   = 8'b00000000; //
            rom[78][1]   = 8'b00000000; //
            rom[78][2]   = 8'b11000110; //**   **
            rom[78][3]   = 8'b11000110; //**   **
            rom[78][4]   = 8'b11100110; //***  **
            rom[78][5]   = 8'b11110110; //**** **
            rom[78][6]   = 8'b11111110; //*******
            rom[78][7]   = 8'b11011110; //** ****
            rom[78][8]   = 8'b11001110; //**  ***
            rom[78][9]   = 8'b11000110; //**   **
            rom[78][10] = 8'b11000110;  //**   **
            rom[78][11] = 8'b11000110;  //**   **
            rom[78][12] = 8'b00000000;  //
            rom[78][13] = 8'b00000000;  //
            rom[78][14] = 8'b00000000;  //
            rom[78][15] = 8'b00000000;  //
            // code x4f (O)
            rom[79][0]   = 8'b00000000; //
            rom[79][1]   = 8'b00000000; //
            rom[79][2]   = 8'b01111100; // *****
            rom[79][3]   = 8'b11111110; //*******
            rom[79][4]   = 8'b11000110; //**   **
            rom[79][5]   = 8'b11000110; //**   **
            rom[79][6]   = 8'b11000110; //**   **
            rom[79][7]   = 8'b11000110; //**   **
            rom[79][8]   = 8'b11000110; //**   **
            rom[79][9]   = 8'b11000110; //**   **
            rom[79][10] = 8'b11111110;  //*******
            rom[79][11] = 8'b01111100;  // *****
            rom[79][12] = 8'b00000000;  //
            rom[79][13] = 8'b00000000;  //
            rom[79][14] = 8'b00000000;  //
            rom[79][15]= 8'b00000000;   //
            // code x50 (P)
            rom[80][0]   = 8'b00000000; //
            rom[80][1]   = 8'b00000000; //
            rom[80][2]   = 8'b11111100; //******
            rom[80][3]   = 8'b11111110; //*******
            rom[80][4]   = 8'b11000110; //**   **
            rom[80][5]   = 8'b11000110; //**   **
            rom[80][6]   = 8'b11111110; //*******
            rom[80][7]   = 8'b11111100; //******   
            rom[80][8]   = 8'b11000000; //**   
            rom[80][9]   = 8'b11000000; //**   
            rom[80][10] = 8'b11000000;  //**
            rom[80][11] = 8'b11000000;  //**
            rom[80][12] = 8'b00000000;  //
            rom[80][13] = 8'b00000000;  //
            rom[80][14] = 8'b00000000;  //
            rom[80][15] = 8'b00000000;  //
            // code x51 (Q)
            rom[81][0]   = 8'b00000000; //
            rom[81][1]   = 8'b00000000; //
            rom[81][2]   = 8'b11111100; // *****
            rom[81][3]   = 8'b11111110; //*******
            rom[81][4]   = 8'b11000110; //**   **
            rom[81][5]   = 8'b11000110; //**   **
            rom[81][6]   = 8'b11000110; //**   **
            rom[81][7]   = 8'b11000110; //**   **  
            rom[81][8]   = 8'b11010110; //** * **
            rom[81][9]   = 8'b11111110; //*******
            rom[81][10] = 8'b01101100;  // ** ** 
            rom[81][11] = 8'b00000110;  //     **
            rom[81][12] = 8'b00000000;  //
            rom[81][13] = 8'b00000000;  //
            rom[81][14] = 8'b00000000;  //
            rom[81][15] = 8'b00000000;  //
            // code x52 (R)
            rom[82][0]   = 8'b00000000; //
            rom[82][1]   = 8'b00000000; //
            rom[82][2]   = 8'b11111100; //******
            rom[82][3]   = 8'b11111110; //*******
            rom[82][4]   = 8'b11000110; //**   **
            rom[82][5]   = 8'b11000110; //**   **
            rom[82][6]   = 8'b11111110; //*******
            rom[82][7]   = 8'b11111100; //******   
            rom[82][8]   = 8'b11011000; //** **  
            rom[82][9]   = 8'b11001100; //**  ** 
            rom[82][10] = 8'b11000110;  //**   **
            rom[82][11] = 8'b11000110;  //**   **
            rom[82][12] = 8'b00000000;  //
            rom[82][13] = 8'b00000000;  //
            rom[82][14] = 8'b00000000;  //
            rom[82][15] = 8'b00000000;  //
            // code x53 (S)
            rom[83][0]   = 8'b00000000; //
            rom[83][1]   = 8'b00000000; //
            rom[83][2]   = 8'b01111100; // *****
            rom[83][3]   = 8'b11111110; //*******
            rom[83][4]   = 8'b11000000; //**   
            rom[83][5]   = 8'b11000000; //**   
            rom[83][6]   = 8'b11111100; //******
            rom[83][7]   = 8'b01111110; // ******   
            rom[83][8]   = 8'b00000110; //     **  
            rom[83][9]   = 8'b00000110; //     **
            rom[83][10] = 8'b11111110;  //*******  
            rom[83][11] = 8'b01111100;  // ***** 
            rom[83][12] = 8'b00000000;  //
            rom[83][13] = 8'b00000000;  //
            rom[83][14] = 8'b00000000;  //
            rom[83][15] = 8'b00000000;  //
            // code x54 (T)
            rom[84][0]   = 8'b00000000; //
            rom[84][1]   = 8'b00000000; //
            rom[84][2]   = 8'b11111110; //*******
            rom[84][3]   = 8'b11111110; //*******
            rom[84][4]   = 8'b00110000; //  **
            rom[84][5]   = 8'b00110000; //  **
            rom[84][6]   = 8'b00110000; //  **
            rom[84][7]   = 8'b00110000; //  **   
            rom[84][8]   = 8'b00110000; //  **  
            rom[84][9]   = 8'b00110000; //  **
            rom[84][10] = 8'b00110000;  //  **  
            rom[84][11] = 8'b00110000;  //  **
            rom[84][12]= 8'b00000000;   //
            rom[84][13] = 8'b00000000;  //
            rom[84][14] = 8'b00000000;  //
            rom[84][15]= 8'b00000000;   //
            // code x55 (U)
            rom[85][0]   = 8'b00000000; //
            rom[85][1]   = 8'b00000000; //
            rom[85][2]   = 8'b11000110; //**   **
            rom[85][3]   = 8'b11000110; //**   **
            rom[85][4]   = 8'b11000110; //**   **
            rom[85][5]   = 8'b11000110; //**   **
            rom[85][6]   = 8'b11000110; //**   **
            rom[85][7]   = 8'b11000110; //**   **
            rom[85][8]   = 8'b11000110; //**   **
            rom[85][9]   = 8'b11000110; //**   **
            rom[85][10] = 8'b11111110;  //*******
            rom[85][11] = 8'b01111100;  // *****
            rom[85][12] = 8'b00000000;  //
            rom[85][13] = 8'b00000000;  //
            rom[85][14] = 8'b00000000;  //
            rom[85][15]= 8'b00000000;   //
            // code x56 (V)
            rom[86][0]   = 8'b00000000; //
            rom[86][1]   = 8'b00000000; //
            rom[86][2]   = 8'b11000110; //**   **
            rom[86][3]   = 8'b11000110; //**   **
            rom[86][4]   = 8'b11000110; //**   **
            rom[86][5]   = 8'b11000110; //**   **
            rom[86][6]   = 8'b11000110; //**   **
            rom[86][7]   = 8'b11000110; //**   **
            rom[86][8]   = 8'b11000110; //**   **
            rom[86][9]   = 8'b01101100; // ** **
            rom[86][10] = 8'b00111000;  //  ***  
            rom[86][11] = 8'b00010000;  //   * 
            rom[86][12] = 8'b00000000;  //
            rom[86][13] = 8'b00000000;  //
            rom[86][14] = 8'b00000000;  //
            rom[86][15]= 8'b00000000;   //
            // code x57 (W)
            rom[87][0]   = 8'b00000000; //
            rom[87][1]   = 8'b00000000; //
            rom[87][2]   = 8'b11000110; //**   **
            rom[87][3]   = 8'b11000110; //**   **
            rom[87][4]   = 8'b11000110; //**   **
            rom[87][5]   = 8'b11000110; //**   **
            rom[87][6]   = 8'b11000110; //**   **
            rom[87][7]   = 8'b11000110; //**   **
            rom[87][8]   = 8'b11010110; //** * **
            rom[87][9]   = 8'b11111110; //*******
            rom[87][10] = 8'b11101110;  //*** ***  
            rom[87][11] = 8'b11000110;  //**   **
            rom[87][12] = 8'b00000000;  //
            rom[87][13] = 8'b00000000;  //
            rom[87][14] = 8'b00000000;  //
            rom[87][15]= 8'b00000000;   //
            // code x58 (X)
            rom[88][0]   = 8'b00000000; //
            rom[88][1]   = 8'b00000000; //
            rom[88][2]   = 8'b11000110; //**   **
            rom[88][3]   = 8'b11000110; //**   **
            rom[88][4]   = 8'b01101100; // ** ** 
            rom[88][5]   = 8'b00111000; //  ***
            rom[88][6]   = 8'b00111000; //  *** 
            rom[88][7]   = 8'b00111000; //  ***
            rom[88][8]   = 8'b00111000; //  ***
            rom[88][9]   = 8'b01101100; // ** **
            rom[88][10] = 8'b11000110;  //**   **  
            rom[88][11] = 8'b11000110;  //**   **
            rom[88][12] = 8'b00000000;  //
            rom[88][13] = 8'b00000000;  //
            rom[88][14] = 8'b00000000;  //
            rom[88][15]= 8'b00000000;   //
            // code x59 (Y)
            rom[89][0]   = 8'b00000000; //
            rom[89][1]   = 8'b00000000; //
            rom[89][2]   = 8'b11000110; //**   **
            rom[89][3]   = 8'b11000110; //**   **
            rom[89][4]   = 8'b01101100; // ** ** 
            rom[89][5]   = 8'b00111000; //  ***
            rom[89][6]   = 8'b00011000; //   ** 
            rom[89][7]   = 8'b00011000; //   **
            rom[89][8]   = 8'b00011000; //   **
            rom[89][9]   = 8'b00011000; //   **
            rom[89][10] = 8'b00011000;  //   **  
            rom[89][11] = 8'b00011000;  //   **
            rom[89][12] = 8'b00000000;  //
            rom[89][13] = 8'b00000000;  //
            rom[89][14] = 8'b00000000;  //
            rom[89][15]= 8'b00000000;   //
            // code x5a (Z)
            rom[90][0]   = 8'b00000000; //
            rom[90][1]   = 8'b00000000; //
            rom[90][2]   = 8'b11111110; //*******
            rom[90][3]   = 8'b11111110; //*******
            rom[90][4]   = 8'b00000110; //     **  
            rom[90][5]   = 8'b00001100; //    **
            rom[90][6]   = 8'b00011000; //   ** 
            rom[90][7]   = 8'b00110000; //  **
            rom[90][8]   = 8'b01100000; // **
            rom[90][9]   = 8'b11000000; //**
            rom[90][10] = 8'b11111110;  //*******  
            rom[90][11] = 8'b11111110;  //*******
            rom[90][12] = 8'b00000000;  //
            rom[90][13] = 8'b00000000;  //
            rom[90][14] = 8'b00000000;  //
            rom[90][15] = 8'b00000000;  //
    end

    always @(*) begin
        pixels = rom[ascii_code][row]; // Output the selected row of the ASCII character
    end

endmodule
